/*----------------------------------------------------------------------------
--     Name    : Note for freq.
--     Made by : Maduinos
--     Date    : 2023/08/19
--     Blog    : https://maduinos.blogspot.com/
--     Ver.    : 0.01
--     WORK    : 
----------------------------------------------------------------------------*/
`define REF_CLK  10000000   // 10Mhz

`define NOTE_B0  (`REF_CLK)/31
`define NOTE_C1  (`REF_CLK)/33
`define NOTE_CS1 (`REF_CLK)/35
`define NOTE_D1  (`REF_CLK)/37
`define NOTE_DS1 (`REF_CLK)/39
`define NOTE_E1  (`REF_CLK)/41
`define NOTE_F1  (`REF_CLK)/44
`define NOTE_FS1 (`REF_CLK)/46
`define NOTE_G1  (`REF_CLK)/49
`define NOTE_GS1 (`REF_CLK)/52
`define NOTE_A1  (`REF_CLK)/55
`define NOTE_AS1 (`REF_CLK)/58
`define NOTE_B1  (`REF_CLK)/62
`define NOTE_C2  (`REF_CLK)/65
`define NOTE_CS2 (`REF_CLK)/69
`define NOTE_D2  (`REF_CLK)/73
`define NOTE_DS2 (`REF_CLK)/78
`define NOTE_E2  (`REF_CLK)/82
`define NOTE_F2  (`REF_CLK)/87
`define NOTE_FS2 (`REF_CLK)/93
`define NOTE_G2  (`REF_CLK)/98
`define NOTE_GS2 (`REF_CLK)/104
`define NOTE_A2  (`REF_CLK)/110
`define NOTE_AS2 (`REF_CLK)/117
`define NOTE_B2  (`REF_CLK)/123
`define NOTE_C3  (`REF_CLK)/131
`define NOTE_CS3 (`REF_CLK)/139
`define NOTE_D3  (`REF_CLK)/147
`define NOTE_DS3 (`REF_CLK)/156
`define NOTE_E3  (`REF_CLK)/165
`define NOTE_F3  (`REF_CLK)/175
`define NOTE_FS3 (`REF_CLK)/185
`define NOTE_G3  (`REF_CLK)/196
`define NOTE_GS3 (`REF_CLK)/208
`define NOTE_A3  (`REF_CLK)/220
`define NOTE_AS3 (`REF_CLK)/233
`define NOTE_B3  (`REF_CLK)/247
`define NOTE_C4  (`REF_CLK)/262
`define NOTE_CS4 (`REF_CLK)/277
`define NOTE_D4  (`REF_CLK)/294
`define NOTE_DS4 (`REF_CLK)/311
`define NOTE_E4  (`REF_CLK)/330
`define NOTE_F4  (`REF_CLK)/349
`define NOTE_FS4 (`REF_CLK)/370
`define NOTE_G4  (`REF_CLK)/392
`define NOTE_GS4 (`REF_CLK)/415
`define NOTE_A4  (`REF_CLK)/440
`define NOTE_AS4 (`REF_CLK)/466
`define NOTE_B4  (`REF_CLK)/494
`define NOTE_C5  (`REF_CLK)/523
`define NOTE_CS5 (`REF_CLK)/554
`define NOTE_D5  (`REF_CLK)/587
`define NOTE_DS5 (`REF_CLK)/622
`define NOTE_E5  (`REF_CLK)/659
`define NOTE_F5  (`REF_CLK)/698
`define NOTE_FS5 (`REF_CLK)/740
`define NOTE_G5  (`REF_CLK)/784
`define NOTE_GS5 (`REF_CLK)/831
`define NOTE_A5  (`REF_CLK)/880
`define NOTE_AS5 (`REF_CLK)/932
`define NOTE_B5  (`REF_CLK)/988
`define NOTE_C6  (`REF_CLK)/1047
`define NOTE_CS6 (`REF_CLK)/1109
`define NOTE_D6  (`REF_CLK)/1175
`define NOTE_DS6 (`REF_CLK)/1245
`define NOTE_E6  (`REF_CLK)/1319
`define NOTE_F6  (`REF_CLK)/1397
`define NOTE_FS6 (`REF_CLK)/1480
`define NOTE_G6  (`REF_CLK)/1568
`define NOTE_GS6 (`REF_CLK)/1661
`define NOTE_A6  (`REF_CLK)/1760
`define NOTE_AS6 (`REF_CLK)/1865
`define NOTE_B6  (`REF_CLK)/1976
`define NOTE_C7  (`REF_CLK)/2093
`define NOTE_CS7 (`REF_CLK)/2217
`define NOTE_D7  (`REF_CLK)/2349
`define NOTE_DS7 (`REF_CLK)/2489
`define NOTE_E7  (`REF_CLK)/2637
`define NOTE_F7  (`REF_CLK)/2794
`define NOTE_FS7 (`REF_CLK)/2960
`define NOTE_G7  (`REF_CLK)/3136
`define NOTE_GS7 (`REF_CLK)/3322
`define NOTE_A7  (`REF_CLK)/3520
`define NOTE_AS7 (`REF_CLK)/3729
`define NOTE_B7  (`REF_CLK)/3951
`define NOTE_C8  (`REF_CLK)/4186
`define NOTE_CS8 (`REF_CLK)/4435
`define NOTE_D8  (`REF_CLK)/4699
`define NOTE_DS8 (`REF_CLK)/4978

